module top_module (
    input clk,
    input d,
    output q
);
    reg q1, q2;
 
    assign q = clk? q1:q2;

    always @ (posedge clk)
        begin
            q1 <= d;
        end

    always @ (negedge clk)
        begin
           q2 <= d; 
        end
    /*
    always @ (posedge clk) begin
    	q1 <= q2^d; 
    end
    
    always @ (negedge clk) begin
    	q2 <= q1^d; 
    end
    //Rising edge，p=d^n, q=d^n^n=d;
    //Falling edge，n=d^p, q=p^d^p=d;
    
    assign q = q1^q2;
    */
endmodule
