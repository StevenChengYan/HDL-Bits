module top_module(
    output zero 
);// Module body starts after semicolon
	zero = 0;
endmodule
